module ej2_gtp2 (
    input wire 
);
    
endmodule